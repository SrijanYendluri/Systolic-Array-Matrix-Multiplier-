`timescale 1ns / 1ps
package mac_uvc_pkg;
	
	`include "uvm_macros.svh"
	import uvm_pkg:: *;
	
	`include "mac_packet.sv" 
	`include "mac_sequence.sv"
	`include "mac_driver.sv"
	`include "mac_monitor.sv"
	`include "mac_agent.sv"
 	`include "mac_scoreboard.sv"
 	`include "env.sv"
// 	`include "mac_top"
	



endpackage